module top_module(
    output zero=0
);
endmodule
